module AND(A,B,O);
  input A;
  input B;
  output O;
  
  and G(O,A,B); //built in AND function
endmodule
